PK   ��S��r�  �    cirkitFile.json��ˎG��w�l[ �����<���@�)����@�|��w�̮[�:l��xc���0�̬�}s=�|~��_���������q��n6?��w������������t�~��>��y�����>�_���Ow�.��L���ͮݽ��]۾:�W���ë��;޼sz�n{���v���n�]���SK3d��.͐U�N�4CVa;�Y��tL3d��m�!����K3d���4CVa;�I3dzF�2-�)@T泲��2-�)�q�����LKt�|d�%:E>4��"�i�N�δD��GgZ����ggZ�S�3-�)��|v��ٙ����LKt�|v�%:E>;��"��i�N��δD��ggZ�w�|v�%:E>;��"��i�Njz>;���LKt�|v�%:E>;��"��i�N��δD��ggZb;�ٙ����LKt�|v�%:E>;��|ș��C>;��"��i�N��δD��ggZ�S�3-�����LKt�|v�%:E>;��"��i�N��δD� _���δD��ggZ�S�3-�)�ٙ��N���LKt�|v�%:E>;W/���������}�a�xy8]�~����{<���k��Y�m��5��k�n;�w;��k�n;�w{��k��w���zG隥��!�wG��k�����zwk��t��m��w�Y�(]�t�������5K���X��X�(]�t�T ~s����k�o�g���v�������k�o�!���a���_��iX���ƹ]�n��a�q�����k�o������a������yX�����t�n��a�q������k�o�	����a�������;�?v�X��������a�q������k�o������a������X����M)����a�q������k�o�NÇ4p��|�{u�?�?,_�|�F ����0߸ˈ�ӧ��1+�?���q��|����?�?,_�|��+����0߸�������5�7nc�p��|�{��?�?,_�|ㆷ�����k�o�M����a�����X����� ��X���Ɠ�������������a�������a�������a�������a������a�������0�x�����0�x2����0�x�����0�x����0�x��O�6���q�8��q����5�7�������5�7�z������5�7�ׅ�����5�7�4f������5�7��������5�7��������g�1����p����6��>����v������z��3DH�y��!��?C���G�z��3DH�y��!���?C���� ��QD��v��r���VJ� bb��Xx+�y`1��n,���<>��X�7�Ji&DL,�w,Ǖ�<Z����o������R�����q�4O"&��;��Ji�EDL,�w,Ǖ�<���8��=�q�4�)"&�I��(�����R����=�q�4�2"&��{��JilDL,�,Ǖ�<战X�X�+�y�1���݇�,�,Ǖ�<	��X�X�+�y.1�?�WJ�$������R�g&��#�q�4OP"&���z�����R��*��#�q�4Y"&��,Ǖ�<r��X�߲���??X��W}>%T�s�\����1�*���u��ixyn��B_+X�k�Ɓ����*���u��ixyψ�B_+X�+�Ɓ����*���u��ixy/��B_+X��Ɓ����*���u��ixy���B_+X׫�Ɓ����*���u��������&z_S�Jh��P/+�-�]5�k5��e��5ի�6���ۚ�UB�zY�mM+�FJ���������^Vz[S�Jh�qS/+���c%��𩗕��T��`��JokjY	m0��e�75���6S���ۚ^VB�zY�m�Wb5�l5r�e��5���6h���ۚ^VB��zY�mM/+��]����������^Vz[��Jh�AX/+���e%��X��������`H��ʓI5���6����ۚ^VB�zY�mM/+��i�����bM/[�zY�mM/+�Fm����������^Vz[��Jh�1\/+���e%��P��������`D��JokzY	m0��e�͆�^VB��zY�mM/+��y����������^Vz[��Jh�A_/+�-�JV��Vc�^Vz[��Jh�!`/+���e%��H��������`@��JokzY	m0.�e��5���6���ftM/+�F�����������^Vz[��Jh�1c/+���e%��б�������`��Jo��Q��V�^Vz[��Jh��d/+���e%�����������`t��JokzY	m0��e哕jzY	m0��e��5���6r���ۚ^�uڿF�?=���`������zz���F���<�L���<�L���<�L���<�L���<�L���<�L���<�L���<�L���<�L���2�l"ҥ��m�ۍ�RZF�����[)-#φ��wc����g��2��WJ�ȳab9�c9����g����7�,�w,Ǖ�2�l�X��X�+�e��0�߱WJ�ȳab9�c9����gS�Y��Y�+�e��0�OR�G),��,Ǖ�2�l�X��Y�+�e��0�߳WJ�ȳab9~`9����g��r��r\)-#φ�}&�>g9~`9����g��r��r\)-#φ�����RZF��W?,Ǐ,Ǖ�2�l�X�Y�+�e��0�o7�כ,Ǐ,Ǖ�2�l�X�Y�+�e��0��e9����g��r����ה��i��i>�:���ȳVe��ȳV��V�#�ā�)>�
}�`F����UZ�Z��<V���*���5y&�nTiU�kk0�LXݦҪ��
�`�8��I�U�����3q`u�J�B_+X��g����V��V�#��|M�Z�&���5���6y��ۢ�Uӻֳ�\Vz[S�Jh��g.+���_%���3����T��h��JokjX	m4��e��5U��6y��ۚ:VB�<sY�mM%+��F���������F#�\V~�P��Jh��g.+���e%���3���}%V��ֳ�\Vz[��Jh��g.+���e%���3�������h��JokzY	m4��e��5���6y��ۚ^VB�<sY�mM/+��F���<�T��Jh��g.+���e%���3�������h��Jo��+����l2�������h��JokzY	m4��e��5���6y��ۚ^VB�<sY�mM/+��F���������F#�\V�l��e%���3�������h��JokzY	m4��e��5���6y��ۢ�d5�l=��e��5���6y��ۚ^VB�<sY�mM/+��F���������F#�\Vz[��Jh��g.+oF����h��JokzY	m4��e��5���6y��ۚ^VB�<sY�mM/+��F������15�l=��e��5���6y��ۚ^VB�<sY�mM/+��F���������F#�\V>Y�����F#�\Vz[��Jh��g.+���e_�����O�����:����y����r=�>>�ޟ����r�;_7o�����t=���s����]��N׻���NG���ˇ�K�ҟ�������7߶'������i�y=:I�����i�y%:I������i�y:I�����i�y�9I������i�e�9["=E|��l @��rs�dh!��X�� GҼƲĜ� Y�@��5���,���ӼƲ����G�R��;��y�e59��t�4���#g9@��@��5��,���ӼƲv��� O� O�˪q�C4|Q�A��A��5���,��=�ӼƲL�� y�y��X�� O O���p����i^cY�r��LŇ� O O��Zp����i^cY�r�<=�<�k,�ُ�A�A��5���,��#�ӼƲ���B���@�A��5���,��#�ӼƲț� yz�4��,�f9@�ނ<]k��.��TNo>���Vu���t�������׻:���/��M���u�G��|�n�����8=���n��wu����,_�k�|���#N��g������]]qz�?���&_��
��#�Y�`�6�zW�<�������������[��xu��Ѳ,4��{�z�
u���R,4�:�	�EX(h<ԕF˯P�x�k	&�^���PWL-�BA㡮'�0Zl���C]Q0a��
����`�h�
�O�uO����*4Ꞃ	�EU(h<�_�螲�"���C�S0a��
����`�h	
uO����)4Ꞃ	�eS(h<�=F�P�x�{
&��J���P�L-�BAs"D�L-�BA��)�0Z���C�S0a�$
���x��)�N(h<�=FˠP�x�{
&�@���P�L-}BA��)�0Z��C�S0a��	����`�h�
��׺�`�h�
uO����&4Ꞃ	�eM(h<�=F�P�xȯ�螲ޞ���C�S0a��	����`�h�
uO����%4Ꞃ	�%K(h<�=F��P��p�=F˔P�x�{
&�(���P�L-MBA��)�0Z����C�S0a�	���ڼ�)��E(h<�=FK�P�x�{
&����P�L-;BA��)�0Zp���I"��`�h�
uO���"#4��q�y�������i��{��o����W>�?�x~���T��g��`�����a�ͧ���G�?~�L����~� o��n�����k?=�?<m~��H���?���tz~U�PK
   ��S��r�  �                  cirkitFile.jsonPK      =   �    